module top_module( input in, output out );
    assign out = !in; // instead of this (!) symbol we can also use (~) this symbol : bitwise negation operator
endmodule
